`include "gate.v"

module main;
reg a, b;
wire abNand, aNot, abAnd, abOr, abXor;

Not  g1(a, aNot);
Nand g2(a, b, aNandb);
And  g3(a, b, aAndb);
Or   g4(a, b, aOrb);
Xor  g5(a, b, aXorb);

initial

begin

  $monitor("%4dns a=%d b=%d aNot=%d abNand=%d abAnd=%d abOr=%d abXor=%d", $stime, a, b, aNot, aNandb, aAndb, aOrb, aXorb);
  a  = 0;
  b  = 0;

end

always #50 begin

  a = a+1;

end

always #100 begin

  b = b+1;

end

initial #500 $finish;

endmodule
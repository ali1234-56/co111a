module hello ;

    initial

        $display ("hello");

endmodule